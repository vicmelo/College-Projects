-------------------------------------------------------------------------
-- Register Bank (R0..R31) - 31 GENERAL PURPOSE 16-bit REGISTERS
-------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_UNSIGNED.all;
use work.p_MR2.all;

entity reg_bank is
	port
	(
		ck, rst, wreg: in std_logic;
		AdRs, AdRt, adRD: in std_logic_vector(4 downto 0);
		RD: in reg32;
		R1, R2: out reg32
	);
end reg_bank;

architecture reg_bank of reg_bank is
	type bank is array(0 to 31) of reg32;
	signal reg: bank;
	signal wen: reg32;
begin

	l1: for i in 0 to 31 generate
		wen(i) <= '1' when i/=0 and adRD=i and wreg='1' else '0';
		-- Remember register $0 is the constant 0, not a register.
		-- This is implemented by never enabling writes to register $0
	end generate l1;
	l2: for i in 0 to 28 generate
		rx: entity work.regnbit generic map(N => 32) port map(ck => ck, rst => rst, ce => wen(i), D => RD, Q => reg(i));
	end generate l2;
	--
	--  Beware! Some registers have specific start values - dependent
	-- on code generation. This version is adapted to work with code
	-- generated by the SPIM simulator
	--
	-- SP ---  x10010000 + x800 -- top of stack
	r29: entity work.regnbit generic map(N => 32, INIT_VALUE => x"10010800") port map(ck => ck, rst => rst, ce => wen(29), D => RD, Q => reg(29));
	r30: entity work.regnbit generic map(N => 32) port map(ck => ck, rst => rst, ce => wen(30), D => RD, Q => reg(30));
	-- $ra --
	r31: entity work.regnbit generic map(N => 32) port map(ck => ck, rst => rst, ce => wen(31), D => RD, Q => reg(31));
	R1 <= reg(CONV_INTEGER(AdRs));	-- source1 selection
	R2 <= reg(CONV_INTEGER(AdRt));	-- source2 selection

end reg_bank;